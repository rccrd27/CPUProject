module multiplier
(
  input [15:0] rs,
  input [15:0] rd,
  output [15:0] q
);

 assign q = ({16{rd[0]}} & {rs[15:0]}) +
				({16{rd[1]}} & {rs[14:0], 1'b0}) +
				({16{rd[2]}} & {rs[13:0], 2'b00}) +
				({16{rd[3]}} & {rs[12:0], 3'b000}) +
				({16{rd[4]}} & {rs[11:0], 4'h0}) +
				({16{rd[5]}} & {rs[10:0], 5'b00000}) +
				({16{rd[6]}} & {rs[9:0], 6'b000000}) +
				({16{rd[7]}} & {rs[8:0], 7'b0000000}) +
				({16{rd[8]}} & {rs[7:0], 8'h00}) +
				({16{rd[9]}} & {rs[6:0], 9'b000000000}) +
				({16{rd[10]}} & {rs[5:0], 10'b0000000000}) +
				({16{rd[11]}} & {rs[4:0], 11'b00000000000}) +
				({16{rd[12]}} & {rs[3:0], 12'h000}) +
				({16{rd[13]}} & {rs[2:0], 13'b0000000000000}) +
				({16{rd[14]}} & {rs[1:0], 14'b00000000000000}) +
				({16{rd[015]}} & {rs[0], 15'b000000000000000});

endmodule 