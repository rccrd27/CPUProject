module Decoder
(
	input [2:0] state,
	input [3:0] inst,
	input [2:0] jmp_flags,
	output [2:0] data_ctrl,
	output e,
	output mux1,
	output WrEn,
	output pc_load,
	output pc_inc,
	output p
	
);
	wire acc_load, mux3, alu;
	wire eq_bar, mi, skip;
	wire lda, sta, add, sub,  jmp, jeq, jmi, stp, ldi, arm;
	wire fetch, exec1, exec2;
	
	assign eq_bar = jmp_flags[2];
	assign mi = jmp_flags[1];
	assign skip = jmp_flags[0];
	
	assign ldi = ~inst[3] & ~inst[2] & ~inst[1] & ~inst[0];
	assign sta = ~inst[3] & ~inst[2] & ~inst[1] & inst[0];
	assign add = ~inst[3] & ~inst[2] & inst[1] & ~inst[0];
	assign sub = ~inst[3] & ~inst[2] & inst[1] & inst[0];
	assign jmp = ~inst[3] & inst[2] & ~inst[1] & ~inst[0];
	assign jmi = ~inst[3] & inst[2] & ~inst[1] & inst[0];
	assign jeq = ~inst[3] & inst[2] & inst[1] & ~inst[0];
	assign stp = ~inst[3] & inst[2] & inst[1] & inst[0];
	assign lda = inst[3] & ~inst[2] & ~inst[1] & ~inst[0];
	assign arm = inst[3] & inst[2];
	
	assign fetch = state[0];
	assign exec1 = state[1];
	assign exec2 = state[2];
	
	assign p = ~fetch & (lda | ldi | jmp | jmi | jeq);
	assign e = lda | add | sub;
	assign mux1 = (exec1 & (lda | jmp | (jmi & mi) | (jeq & ~eq_bar))) | (~fetch & (sta | add | sub));
	assign WrEn = exec1 & sta;
	assign pc_load = (exec1 | fetch & skip) & (jmp | (jmi & mi) | (jeq & ~eq_bar));
	assign pc_inc = exec1 & ~(stp | jmp | (jmi & mi) | (jeq & ~eq_bar));
	assign acc_load = (exec1 & ldi) | (exec2 & (lda | add | sub));
	assign mux3 = add | sub;
	assign alu = add;
	
	assign data_ctrl = {alu, mux3, acc_load};

endmodule

