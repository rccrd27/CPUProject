module multiplier
(
  input [15:0] rs,
  input [15:0] rd,
  output [15:0] q
);

 assign q = rd[0] & {rs[15:0]} +
				rd[1] & {rs[14:0], 1'h0} +
				rd[2] & {rs[13:0], 2'h0} +
				rd[3] & {rs[12:0], 3'h0} +
				rd[4] & {rs[11:0], 4'h0} +
				rd[5] & {rs[10:0], 5'h00} +
				rd[6] & {rs[9:0], 6'h00} +
				rd[7] & {rs[8:0], 7'h00} +
				rd[8] & {rs[7:0], 8'h00} +
				rd[9] & {rs[6:0], 9'h000} +
				rd[10] & {rs[5:0], 10'h000} +
				rd[11] & {rs[4:0], 11'h000} +
				rd[12] & {rs[3:0], 12'h000} +
				rd[13] & {rs[2:0], 13'h0000} +
				rd[14] & {rs[1:0], 14'h0000} +
				rd[15] & {rs[0], 15'h0000};

endmodule 